`timescale 1ns/10ps


module cla19(A,B,Cin,Sum);
input[18:0]A,B;
input Cin;
output[18:0]Sum;
//output Cout;
wire G,P;
wire [18:0]B_,gtemp1,ptemp1,ctemp1;
wire [3:0]gouta,pouta;
wire [4:0] ctemp2;
wire t1,t2,t3,t4;
xor(B_[0],B[0],Cin);
xor(B_[1],B[1],Cin);
xor(B_[2],B[2],Cin);
xor(B_[3],B[3],Cin);
xor(B_[4],B[4],Cin);
xor(B_[5],B[5],Cin);
xor(B_[6],B[6],Cin);
xor(B_[7],B[7],Cin);
xor(B_[8],B[8],Cin);
xor(B_[9],B[9],Cin);
xor(B_[10],B[10],Cin);
xor(B_[11],B[11],Cin);
xor(B_[12],B[12],Cin);
xor(B_[13],B[13],Cin);
xor(B_[14],B[14],Cin);
xor(B_[15],B[15],Cin);
xor(B_[16],B[16],Cin);
xor(B_[17],B[17],Cin);
xor(B_[18],B[18],Cin);
RFA r01 (gtemp1[0],ptemp1[0],Sum[0],A[0],B_[0],Cin);
RFA r02 (gtemp1[1],ptemp1[1],Sum[1],A[1],B_[1],ctemp1[1]);
RFA r03 (gtemp1[2],ptemp1[2],Sum[2],A[2],B_[2],ctemp1[2]);
RFA r04 (gtemp1[3],ptemp1[3],Sum[3],A[3],B_[3],ctemp1[3]);
bclg4 b1(ctemp1[3:0],gouta[0],pouta[0],gtemp1[3:0],ptemp1[3:0],Cin);
RFA r05 (gtemp1[4],ptemp1[4],Sum[4],A[4],B_[4],ctemp2[1]);
RFA r06 (gtemp1[5],ptemp1[5],Sum[5],A[5],B_[5],ctemp1[5]);
RFA r07 (gtemp1[6],ptemp1[6],Sum[6],A[6],B_[6],ctemp1[6]);
RFA r08 (gtemp1[7],ptemp1[7],Sum[7],A[7],B_[7],ctemp1[7]);
bclg4 b2(ctemp1[7:4],gouta[1],pouta[1],gtemp1[7:4],ptemp1[7:4],ctemp2[1]);
RFA r09 (gtemp1[8],ptemp1[8],Sum[8],A[8],B_[8],ctemp2[2]);
RFA r10 (gtemp1[9],ptemp1[9],Sum[9],A[9],B_[9],ctemp1[9]);
RFA r11 (gtemp1[10],ptemp1[10],Sum[10],A[10],B_[10],ctemp1[10]);
RFA r12 (gtemp1[11],ptemp1[11],Sum[11],A[11],B_[11],ctemp1[11]);
bclg4 b3(ctemp1[11:8],gouta[2],pouta[2],gtemp1[11:8],ptemp1[11:8],ctemp2[2]);
RFA r13 (gtemp1[12],ptemp1[12],Sum[12],A[12],B_[12],ctemp2[3]);
RFA r14 (gtemp1[13],ptemp1[13],Sum[13],A[13],B_[13],ctemp1[13]);
RFA r15 (gtemp1[14],ptemp1[14],Sum[14],A[14],B_[14],ctemp1[14]);
RFA r16 (gtemp1[15],ptemp1[15],Sum[15],A[15],B_[15],ctemp1[15]);
bclg4 b4(ctemp1[15:12],gouta[3],pouta[3],gtemp1[15:12],ptemp1[15:12],ctemp2[3]);
bclg4 b5(ctemp2[3:0],G,P,gouta,pouta,Cin);
RFA r17 (gtemp1[16],ptemp1[16],Sum[16],A[16],B_[16],ctemp2[4]);
RFA r18 (gtemp1[17],ptemp1[17],Sum[17],A[17],B_[17],ctemp1[17]);
RFA r19 (gtemp1[18],ptemp1[18],Sum[18],A[18],B_[18],ctemp1[18]);
and(t1,P,Cin);
or(ctemp2[4],G,t1);
and(t2,ptemp1[16],ctemp2[4]);
or(ctemp1[17],gtemp1[16],t2);
and(t3,ptemp1[17],gtemp1[16]);
and(t4,ptemp1[17],ptemp1[16],ctemp2[4]);
or(ctemp1[18],gtemp1[17],t3,t4);
/*and(t5,ptemp1[18],ctemp1[17]);
or(Cout,gtemp1[18],t5);*/
endmodule